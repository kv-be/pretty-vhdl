-------------
-- begin
-------------




---------     
-- END
---------
